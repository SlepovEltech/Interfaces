library verilog;
use verilog.vl_types.all;
entity UART_vlg_vec_tst is
end UART_vlg_vec_tst;
