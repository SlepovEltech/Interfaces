library verilog;
use verilog.vl_types.all;
entity sinus_vlg_sample_tst is
    port(
        QUARZ           : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end sinus_vlg_sample_tst;
