library verilog;
use verilog.vl_types.all;
entity sinus_vlg_vec_tst is
end sinus_vlg_vec_tst;
